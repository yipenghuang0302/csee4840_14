`timescale 1ns/1ps
`include "cholesky_test.sv"

class cholesky_transaction;
	rand logic [6][6][30:0] j_increment;
	real j_fraction [6][6];
	real j_data [6][6];
	real matrix_data [6][6];
endclass

class cholesky_env;
	int max_transactions = 1000000;
endclass

program cholesky_tb (ifc_cholesky.cholesky_tb ds);

	cholesky_transaction trans;
	cholesky_env env;
	cholesky_test test;

	task do_cycle;

		trans.randomize();

		//wrap input numbers to -16 ~ 16
		for ( int row=0 ; row<6 ; row++ ) begin // row index
			for ( int col=0 ; col<6 ; col++ ) begin // col index
				trans.j_fraction[row][col] = real'(trans.j_increment[row][col]) / 2147483648.0;
				trans.j_data[row][col] = -16.0 + trans.j_fraction[row][col] * 2 * 16.0;
			end
		end

		// create jjt which is positive symmetric definite
		for ( int row=0 ; row<6 ; row++ ) begin // row index
			for ( int col=0 ; col<6 ; col++ ) begin // col index
				trans.matrix_data[row][col] = 0.0;
				for ( int index=0 ; index<6 ; index++ ) begin // index
					trans.matrix_data[row][col] += trans.j_data[row][index] * trans.j_data[col][index];
				end
				$display("row, col = %d", row, col);
				$display("data = %f", trans.matrix_data[row][col]);
				ds.cb.matrix[row][col] <= int'(trans.matrix_data[row][col] * 256.0);
			end
		end

		ds.cb.en <= 1'b1;
		ds.cb.rst <= 1'b0;

		@(ds.cb);
		test.update_cholesky (
			trans.matrix_data
		);

	endtask

	initial begin
		trans = new();
		test = new();
		env = new();

		@(ds.cb);
		ds.cb.rst <= 1'b1;
		@(ds.cb);

		// testing
		repeat (env.max_transactions) begin
			do_cycle();
			repeat (210) @(ds.cb);
			test.check_cholesky (
				ds.cb.lt
			);
		end
	end
endprogram