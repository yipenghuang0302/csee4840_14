// megafunction wizard: %ALTSQRT%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: ALTSQRT 

// ============================================================
// File Name: sqrt_27.v
// Megafunction Name(s):
// 			ALTSQRT
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 13.1.3 Build 178 02/12/2014 SJ Web Edition
// ************************************************************


//Copyright (C) 1991-2014 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module sqrt_27 (
	clk,
	ena,
	radical,
	q,
	remainder);

	input	  clk;
	input	  ena;
	input	[26:0]  radical;
	output	[13:0]  q;
	output	[14:0]  remainder;

	wire [13:0] sub_wire0;
	wire [14:0] sub_wire1;
	wire [13:0] q = sub_wire0[13:0];
	wire [14:0] remainder = sub_wire1[14:0];

	altsqrt	ALTSQRT_component (
				.clk (clk),
				.ena (ena),
				.radical (radical),
				.q (sub_wire0),
				.remainder (sub_wire1)
				// synopsys translate_off
				,
				.aclr ()
				// synopsys translate_on
				);
	defparam
		ALTSQRT_component.pipeline = 5,
		ALTSQRT_component.q_port_width = 14,
		ALTSQRT_component.r_port_width = 15,
		ALTSQRT_component.width = 27;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "1"
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: CONSTANT: PIPELINE NUMERIC "5"
// Retrieval info: CONSTANT: Q_PORT_WIDTH NUMERIC "14"
// Retrieval info: CONSTANT: R_PORT_WIDTH NUMERIC "15"
// Retrieval info: CONSTANT: WIDTH NUMERIC "27"
// Retrieval info: USED_PORT: clk 0 0 0 0 INPUT NODEFVAL "clk"
// Retrieval info: USED_PORT: ena 0 0 0 0 INPUT NODEFVAL "ena"
// Retrieval info: USED_PORT: q 0 0 14 0 OUTPUT NODEFVAL "q[13..0]"
// Retrieval info: USED_PORT: radical 0 0 27 0 INPUT NODEFVAL "radical[26..0]"
// Retrieval info: USED_PORT: remainder 0 0 15 0 OUTPUT NODEFVAL "remainder[14..0]"
// Retrieval info: CONNECT: @clk 0 0 0 0 clk 0 0 0 0
// Retrieval info: CONNECT: @ena 0 0 0 0 ena 0 0 0 0
// Retrieval info: CONNECT: @radical 0 0 27 0 radical 0 0 27 0
// Retrieval info: CONNECT: q 0 0 14 0 @q 0 0 14 0
// Retrieval info: CONNECT: remainder 0 0 15 0 @remainder 0 0 15 0
// Retrieval info: GEN_FILE: TYPE_NORMAL sqrt_27.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL sqrt_27.inc TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL sqrt_27.cmp TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL sqrt_27.bsf TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL sqrt_27_inst.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL sqrt_27_bb.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL sqrt_27_syn.v TRUE
// Retrieval info: LIB_FILE: altera_mf
