// megafunction wizard: %ALTSQRT%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: ALTSQRT 

// ============================================================
// File Name: sqrt_43.v
// Megafunction Name(s):
// 			ALTSQRT
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 13.1.4 Build 182 03/12/2014 SJ Web Edition
// ************************************************************


//Copyright (C) 1991-2014 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module sqrt_43 (
	clk,
	ena,
	radical,
	q,
	remainder);

	input	  clk;
	input	  ena;
	input	[42:0]  radical;
	output	[21:0]  q;
	output	[22:0]  remainder;

	wire [21:0] sub_wire0;
	wire [22:0] sub_wire1;
	wire [21:0] q = sub_wire0[21:0];
	wire [22:0] remainder = sub_wire1[22:0];

	altsqrt	ALTSQRT_component (
				.clk (clk),
				.ena (ena),
				.radical (radical),
				.q (sub_wire0),
				.remainder (sub_wire1)
				// synopsys translate_off
				,
				.aclr ()
				// synopsys translate_on
				);
	defparam
		ALTSQRT_component.pipeline = 5,
		ALTSQRT_component.q_port_width = 22,
		ALTSQRT_component.r_port_width = 23,
		ALTSQRT_component.width = 43;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: CONSTANT: PIPELINE NUMERIC "5"
// Retrieval info: CONSTANT: Q_PORT_WIDTH NUMERIC "22"
// Retrieval info: CONSTANT: R_PORT_WIDTH NUMERIC "23"
// Retrieval info: CONSTANT: WIDTH NUMERIC "43"
// Retrieval info: USED_PORT: clk 0 0 0 0 INPUT NODEFVAL "clk"
// Retrieval info: USED_PORT: ena 0 0 0 0 INPUT NODEFVAL "ena"
// Retrieval info: USED_PORT: q 0 0 22 0 OUTPUT NODEFVAL "q[21..0]"
// Retrieval info: USED_PORT: radical 0 0 43 0 INPUT NODEFVAL "radical[42..0]"
// Retrieval info: USED_PORT: remainder 0 0 23 0 OUTPUT NODEFVAL "remainder[22..0]"
// Retrieval info: CONNECT: @clk 0 0 0 0 clk 0 0 0 0
// Retrieval info: CONNECT: @ena 0 0 0 0 ena 0 0 0 0
// Retrieval info: CONNECT: @radical 0 0 43 0 radical 0 0 43 0
// Retrieval info: CONNECT: q 0 0 22 0 @q 0 0 22 0
// Retrieval info: CONNECT: remainder 0 0 23 0 @remainder 0 0 23 0
// Retrieval info: GEN_FILE: TYPE_NORMAL sqrt_43.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL sqrt_43.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL sqrt_43.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL sqrt_43.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL sqrt_43_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL sqrt_43_bb.v FALSE
// Retrieval info: LIB_FILE: altera_mf
