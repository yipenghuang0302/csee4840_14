module divider (input clk, 
                input div_en,
                input [4:0][26:0] dividends, 
                input [26:0] divisor,
                output [4:0][26:0] quotients);

endmodule
